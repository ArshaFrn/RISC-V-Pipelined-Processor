module InstructionMemory(input logic [31:0] addr, 
                         output logic [31:0] instruction);
    logic [31:0] instruction_memory [31:0];    
    initial begin
        $readmemh("E:\\University\\CA\\Project\\RISC-V-Pipelined-Processor\\src\\code2.mem", instruction_memory);
    end
    assign instruction = instruction_memory[addr[31:2]];
endmodule
